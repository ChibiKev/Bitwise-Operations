library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Chen_Kevin_Rotation_Right_tb is
end Chen_Kevin_Rotation_Right_tb;

architecture Chen_Kevin_tb of Chen_Kevin_Rotation_Right_tb is
    signal Chen_Kevin_a: std_logic_vector(5 downto 0);  -- inputs 
    signal Chen_Kevin_result : std_logic_vector(5 downto 0);  -- outputs
begin

    UUT : entity work.Chen_Kevin_Rotation_Right port map (Chen_Kevin_a => Chen_Kevin_a,
																		Chen_Kevin_result => Chen_Kevin_result);
		process
		begin
		
		Chen_Kevin_a <= "000000";
		
		for i in 0 to 63
		loop
		wait for 10 ns;
		Chen_Kevin_a <= std_logic_vector(unsigned(Chen_Kevin_a) + 1);
		end loop;
		
		end process;
end Chen_Kevin_tb;